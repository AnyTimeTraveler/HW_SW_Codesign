-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW(7-0) are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY(0) is the active-low system reset
-- Outputs: LEDG(7-0) are parallel outputs from the Nios system
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY aufgabe4 IS
	PORT(
		KEY      : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
		CLOCK_50 : IN STD_LOGIC
	);
END aufgabe4;

ARCHITECTURE structure OF aufgabe4 IS

	 component nios_system is
		port (
			clk_clk       : in std_logic;
			reset_reset_n : in std_logic
		);
	end component nios_system;

BEGIN
	-- Instantiate the Nios system entity generated by Qsys
	myNios_inst : nios_system
		PORT MAP(
			clk_clk       => CLOCK_50,
			reset_reset_n => KEY(0)
		);

END structure;
