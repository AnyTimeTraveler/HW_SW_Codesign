-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW(7-0) are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY(0) is the active-low system reset
-- Outputs: LEDG(7-0) are parallel outputs from the Nios system
LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY lights IS
PORT (
	SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLOCK_50 : IN STD_LOGIC;
	LEDG : OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
END lights;

ARCHITECTURE structure OF lights IS
COMPONENT nios_system PORT (
	-- 1) global signals:
	clk_clk : IN STD_LOGIC;
	reset_reset_n : IN STD_LOGIC;
	-- the_pio_leds
	pio_leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	-- the_pio_switches
	pio_switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

BEGIN
-- Instantiate the Nios system entity generated by Qsys
myNios_inst : nios_system PORT MAP(
		pio_leds_export => LEDG(7 DOWNTO 0),
		clk_clk => CLOCK_50,
		pio_switches_export => SW(7 DOWNTO 0),
		reset_reset_n => KEY(0) );
END structure;
