-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW(7-0) are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY(0) is the active-low system reset
-- Outputs: LEDG(7-0) are parallel outputs from the Nios system
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY aufgabe3 IS
	PORT(
		SW							   : IN	STD_LOGIC_VECTOR(17 DOWNTO 0);
		KEY							  : IN	STD_LOGIC_VECTOR(3 DOWNTO 0);
		CLOCK_50						 : IN	STD_LOGIC;
		LEDG							 : OUT   STD_LOGIC_VECTOR(8 DOWNTO 0);
		LEDR							 : OUT   STD_LOGIC_VECTOR(7 DOWNTO 0);
		-- SDRAM signals
		DRAM_DQ						  : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
		DRAM_ADDR						: OUT   STD_LOGIC_VECTOR(12 DOWNTO 0);
		DRAM_BA						  : OUT   STD_LOGIC_VECTOR(1 DOWNTO 0);
		DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK : OUT   STD_LOGIC;
		DRAM_CKE, DRAM_CS_N, DRAM_WE_N   : OUT   STD_LOGIC;
		DRAM_DQM						 : OUT   STD_LOGIC_VECTOR(3 DOWNTO 0);
		UART_RXD		   		: in	std_logic					 := 'X';			 -- RXD
		UART_TXD		   		: out   std_logic;										-- TXD
		LCD_RS			  : out   std_logic;										-- RS
		LCD_RW			  : out   std_logic;										-- RW
		LCD_DATA 			: inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
		LCD_EN			   : out   std_logic										 -- E
	);
END aufgabe3;

ARCHITECTURE structure OF aufgabe3 IS
	COMPONENT pll
		PORT(
			inclk0 : in  std_logic;
			c0	 : out std_logic;
			c1	 : out std_logic
		);
	END COMPONENT;

	 component nios_system is
		port (
			clk_clk			 : in	std_logic					 := 'X';			 -- clk
			pio_leds_export	 : out   std_logic_vector(15 downto 0);					-- export
			pio_switches_export : in	std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			reset_reset_n	   : in	std_logic					 := 'X';			 -- reset_n
			sdram_wire_addr	 : out   std_logic_vector(12 downto 0);					-- addr
			sdram_wire_ba	   : out   std_logic_vector(1 downto 0);					 -- ba
			sdram_wire_cas_n	: out   std_logic;										-- cas_n
			sdram_wire_cke	  : out   std_logic;										-- cke
			sdram_wire_cs_n	 : out   std_logic;										-- cs_n
			sdram_wire_dq	   : inout std_logic_vector(31 downto 0) := (others => 'X'); -- dq
			sdram_wire_dqm	  : out   std_logic_vector(3 downto 0);					 -- dqm
			sdram_wire_ras_n	: out   std_logic;										-- ras_n
			sdram_wire_we_n	 : out   std_logic;										-- we_n
			rs232_RXD		   : in	std_logic					 := 'X';			 -- RXD
			rs232_TXD		   : out   std_logic;										-- TXD
			lcd_RS			  : out   std_logic;										-- RS
			lcd_RW			  : out   std_logic;										-- RW
			lcd_data			: inout std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			lcd_E			   : out   std_logic										 -- E
		);
	end component nios_system;


	SIGNAL counter_output : std_ulogic_vector(31 downto 0);
	SIGNAL pio_leds	   : std_logic_vector(15 downto 0);
	SIGNAL cpu_clk		: std_logic;
	SIGNAL sdram_clk	  : std_logic;

BEGIN
	pll_inst : pll
		PORT MAP (
			inclk0 => CLOCK_50,
			c0	 => cpu_clk,
			c1	 => sdram_clk
		);

	-- Instantiate the Nios system entity generated by Qsys
	myNios_inst : nios_system
		PORT MAP(
			clk_clk				=> CLOCK_50,
			pio_leds_export		=> pio_leds,
			pio_switches_export	=> SW(7 downto 0),
			reset_reset_n		=> KEY(0),
			sdram_wire_addr		=> DRAM_ADDR,
			sdram_wire_ba		=> DRAM_BA,
			sdram_wire_cas_n	=> DRAM_CAS_N,
			sdram_wire_cke		=> DRAM_CKE,
			sdram_wire_cs_n		=> DRAM_CS_N,
			sdram_wire_dq		=> DRAM_DQ,
			sdram_wire_dqm		=> DRAM_DQM,
			sdram_wire_ras_n	=> DRAM_RAS_N,
			sdram_wire_we_n		=> DRAM_WE_N,
			rs232_RXD			=> UART_RXD,
			rs232_TXD			=> UART_TXD,
			lcd_RS				=> LCD_RS,
			lcd_RW				=> LCD_RW,
			lcd_data			=> LCD_DATA(7 downto 0),
			lcd_E				=> LCD_EN
		);


	LEDG(7 DOWNTO 0) <= pio_leds(7 downto 0);
	LEDR(7 DOWNTO 0) <= pio_leds(15 downto 8);
	DRAM_CLK		 <= sdram_clk;
END structure;
