-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW(7-0) are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY(0) is the active-low system reset
-- Outputs: LEDG(7-0) are parallel outputs from the Nios system
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY lights IS
PORT (
        SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
        KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
        CLOCK_50 : IN STD_LOGIC;
        LEDG : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        LEDR : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
        -- SDRAM signals
        DRAM_DQ : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
        DRAM_ADDR : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
        DRAM_BA : OUT STD_LOGIC_VECTOR (1 DOWNTO 0);
        DRAM_CAS_N, DRAM_RAS_N, DRAM_CLK : OUT STD_LOGIC;
        DRAM_CKE, DRAM_CS_N, DRAM_WE_N : OUT STD_LOGIC;
        DRAM_DQM : OUT STD_LOGIC_VECTOR (3 DOWNTO 0)
);
END lights;

ARCHITECTURE structure OF lights IS
COMPONENT nios_system PORT (
        clk_clk             : in    std_logic;
        pio_leds_export     : out   std_logic_vector(15 downto 0);
        pio_switches_export : in    std_logic_vector(7 downto 0);
        reset_reset_n       : in    std_logic;
        sdram_wire_addr     : out   std_logic_vector(12 downto 0);
        sdram_wire_ba       : out   std_logic_vector(1 downto 0);
        sdram_wire_cas_n    : out   std_logic;
        sdram_wire_cke      : out   std_logic;
        sdram_wire_cs_n     : out   std_logic;
        sdram_wire_dq       : inout std_logic_vector(31 downto 0);
        sdram_wire_dqm      : out   std_logic_vector(3 downto 0);
        sdram_wire_ras_n    : out   std_logic;
        sdram_wire_we_n     : out   std_logic
);
END COMPONENT;

COMPONENT counter
        GENERIC (
                BIT_WIDTH: integer
        );
        PORT
        (
                clk                 : in std_ulogic;
                reset_n         : in std_ulogic;
                enable         : in std_ulogic;
                q                 : out std_ulogic_vector(BIT_WIDTH - 1 downto 0)
        );

END COMPONENT;

SIGNAL counter_output : std_ulogic_vector(31 downto 0);
SIGNAL pio_leds : std_logic_vector(15 downto 0);

BEGIN
-- Instantiate the Nios system entity generated by Qsys
myNios_inst : nios_system PORT MAP(
        clk_clk => CLOCK_50,
        pio_leds_export => pio_leds,
        pio_switches_export => SW(7 downto 0),
        reset_reset_n => KEY(0),
        sdram_wire_addr => DRAM_ADDR,
        sdram_wire_ba => DRAM_BA,
        sdram_wire_cas_n => DRAM_CAS_N,
        sdram_wire_cke => DRAM_CKE,
        sdram_wire_cs_n => DRAM_CS_N,
        sdram_wire_dq => DRAM_DQ,
        sdram_wire_dqm => DRAM_DQM,
        sdram_wire_ras_n => DRAM_RAS_N,
        sdram_wire_we_n => DRAM_WE_N
);

counter_inst: counter
        GENERIC MAP(
                BIT_WIDTH => 32
        )
        PORT MAP
        (
                clk                 => CLOCK_50,
                reset_n         => KEY(0),
                enable         => '1',
                q                  => counter_output
        );
        
process(counter_output, pio_leds)
        variable offset : unsigned(7 downto 0);
begin
        offset := unsigned(pio_leds(7 downto 0));
        LEDG(8) <= counter_output(20 + to_integer(offset));
end process;

LEDG(7 DOWNTO 0) <= pio_leds(7 downto 0);
LEDR(7 DOWNTO 0) <= pio_leds(15 downto 8);
DRAM_CLK <= CLOCK_50;
END structure;