-- Implements a simple Nios II system for the DE2-115 board.
-- Inputs: SW(7-0) are parallel port inputs to the Nios II system
-- CLOCK_50 is the system clock
-- KEY(0) is the active-low system reset
-- Outputs: LEDG(7-0) are parallel outputs from the Nios system
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use ieee.numeric_std.all;

ENTITY lights IS
PORT (
	SW : IN STD_LOGIC_VECTOR(17 DOWNTO 0);
	KEY : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
	CLOCK_50 : IN STD_LOGIC;
	LEDG : OUT STD_LOGIC_VECTOR(8 DOWNTO 0));
END lights;

ARCHITECTURE structure OF lights IS
COMPONENT nios_system PORT (
	-- 1) global signals:
	clk_clk : IN STD_LOGIC;
	reset_reset_n : IN STD_LOGIC;
	-- the_pio_leds
	pio_leds_export : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	-- the_pio_switches
	pio_switches_export : IN STD_LOGIC_VECTOR(7 DOWNTO 0));
END COMPONENT;

COMPONENT counter
	GENERIC (
		BIT_WIDTH: integer
	);
	PORT
	(
		clk		 : in std_ulogic;
		reset_n	 : in std_ulogic;
		enable	 : in std_ulogic;
		q		 : out std_ulogic_vector(BIT_WIDTH - 1 downto 0)
	);

END COMPONENT;

SIGNAL counter_output : std_ulogic_vector(31 downto 0);
SIGNAL pio_leds : std_logic_vector(7 downto 0);

BEGIN
-- Instantiate the Nios system entity generated by Qsys
myNios_inst : nios_system PORT MAP(
		pio_leds_export => pio_leds,
		clk_clk => CLOCK_50,
		pio_switches_export => SW(7 DOWNTO 0),
		reset_reset_n => KEY(0) );
		
counter_inst: counter
	GENERIC MAP(
		BIT_WIDTH => 32
	)
	PORT MAP
	(
		clk		 => CLOCK_50,
		reset_n	 => KEY(0),
		enable	 => '1',
		q		  => counter_output
	);
	
process(counter_output, pio_leds)
	variable offset : unsigned(7 downto 0);
begin
	offset := unsigned(pio_leds);
	LEDG(8) <= counter_output(20 + to_integer(offset));
end process;
	
LEDG(7 DOWNTO 0) <= pio_leds;
END structure;
